module I2S_Slave(clk, rst_n, I2S_sclk, I2S_ws, I2S_data,
		 lft_chnnl, rght_chnnl, vld);

input clk, rst_n, I2S_sclk, I2S_ws, I2S_data;
output [23:0] lft_chnnl, rght_chnnl;
output reg vld;

//////////////////////
// sclk rise detect //
//////////////////////
wire sclk_rise;
reg sclk_FF1, sclk_FF2, sclk_FF3;
// Double flop for metastability
always_ff @ (posedge clk, negedge rst_n)
	if(!rst_n) begin
		sclk_FF1 <= 1'b0;
		sclk_FF2 <= 1'b0;
		sclk_FF3 <= 1'b0;
	end
	else begin
		sclk_FF1 <= I2S_sclk;
		sclk_FF2 <= sclk_FF1;
		sclk_FF3 <= sclk_FF2;
	end
assign sclk_rise = ~sclk_FF3 & sclk_FF2;

////////////////////
// ws_fall detect //
////////////////////
wire ws_fall;
reg ws_FF1, ws_FF2, ws_FF3;
// Double flop for metastability
always_ff @ (posedge clk, negedge rst_n)
	if(!rst_n) begin
		ws_FF1 <= 1'b0;
		ws_FF2 <= 1'b0;
		ws_FF3 <= 1'b0;
	end
	else begin
		ws_FF1 <= I2S_ws;
		ws_FF2 <= ws_FF1;
		ws_FF3 <= ws_FF2;
	end
assign ws_fall = ws_FF3 & ~ws_FF2;

////////////////////
// Shift register //
////////////////////
reg[47:0] shft_reg;
always @ (posedge clk, negedge rst_n)
	if(!rst_n) shft_reg <= 48'd0;
	else if(sclk_rise) shft_reg <= {shft_reg[46:0], I2S_data};

assign lft_chnnl = shft_reg[47:24];
assign rght_chnnl = shft_reg[23:0];

/////////////
// Counter //
/////////////
reg[4:0] bit_cntr;
reg clr_cnt;
wire eq22, eq24;

always @ (posedge clk, negedge rst_n)
	if(!rst_n) bit_cntr <= 5'h00;
	else if(clr_cnt) bit_cntr <= 5'h00;
	else if(sclk_rise) bit_cntr <= bit_cntr + 1'b1;
assign eq22 = (bit_cntr == 5'd22) ? 1'b1 : 1'b0;
assign eq24 = (bit_cntr == 5'd24) ? 1'b1 : 1'b0;

///////////////////
// State machine //
///////////////////
typedef enum reg[1:0] {SYNC, SKIP, LEFT, RIGHT} state_t;
state_t state, nxt;

reg set_val;

always_ff @ (posedge clk, negedge rst_n)
	if(!rst_n) state <= SYNC;
	else state <= nxt;

always_comb begin
	clr_cnt = 0;
	set_val = 0;
	nxt = SYNC;

	case(state)
	 SYNC: 
		if(ws_fall) nxt = SKIP;
	 SKIP: 
		if(sclk_rise) begin 
			nxt = LEFT;
			clr_cnt = 1;
		end
		else nxt = SKIP;
	 LEFT:
		if(eq24) begin	
			nxt = RIGHT;
			clr_cnt = 1;
		end
		else nxt = LEFT;
	RIGHT:
		if(eq24) begin
			nxt = LEFT;
			clr_cnt = 1;
			set_val = 1;
		end
		else if(eq22 & !I2S_ws)
			nxt = SYNC;
		else nxt = RIGHT;
	endcase
end

///////////////////////////////
// Set valid (one clk cycle) //
///////////////////////////////
always @ (posedge clk, negedge rst_n)
	if(!rst_n) vld <= 1'b0;
	else vld <= set_val;

endmodule 
