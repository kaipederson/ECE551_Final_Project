module LED();

endmodule
